
`timescale 1 ns / 1 ps

	module systolic_array #
	(
		// Users to add parameters here
	parameter SYSTOLIC_SIZE     = 16      ,
	parameter DATA_WIDTH        = 16      ,
	parameter INOUT_WIDTH       = 256     ,
	parameter IFM_RAM_SIZE      = 524172  ,
	parameter WGT_RAM_SIZE      = 5040 ,
	parameter OFM_RAM_SIZE_1    = 2205619 ,
  parameter OFM_RAM_SIZE_2    = 259584  ,
	parameter MAX_WGT_FIFO_SIZE = 4608    ,
	parameter RELU_PARAM        = 0       ,
  parameter Q                 = 9       ,
  parameter NUM_LAYER         = 1       ,
  parameter ID_WIDTH          = 4       ,
  parameter ADDR_WIDTH        = 32      ,
  parameter LEN_WIDTH         = 8       ,


		// Parameters of Axi Master Bus Interface M00_AXI

		parameter  C_M_TARGET_SLAVE_BASE_ADDR  = 32'h40000000,
		parameter integer C_M_AXI_BURST_LEN    = 256,
		parameter integer C_M_AXI_ID_WIDTH     = 4,
		parameter integer C_M_AXI_ADDR_WIDTH   = 32,
		parameter integer C_M_AXI_DATA_WIDTH   = 256,
		parameter integer C_M_AXI_AWUSER_WIDTH = 0,
		parameter integer C_M_AXI_ARUSER_WIDTH = 0,
		parameter integer C_M_AXI_WUSER_WIDTH  = 0,
		parameter integer C_M_AXI_RUSER_WIDTH  = 0,
		parameter integer C_M_AXI_BUSER_WIDTH  = 0

	)
	(
		// Users to add ports here

		// User ports ends
		// Do not modify the ports beyond this line


		// Ports of Axi Master Bus Interface M00_AXI
		input wire                                 m00_axi_init_axi_txn ,
		output wire                                m00_axi_txn_done     ,
		output wire                                m00_axi_error        ,
		input wire                                 m00_axi_aclk         ,
		input wire                                 m00_axi_aresetn      ,
		output wire [C_M00_AXI_ID_WIDTH-1 : 0]     m00_axi_awid         ,
		output wire [C_M00_AXI_ADDR_WIDTH-1 : 0]   m00_axi_awaddr       ,
		output wire [7 : 0]                        m00_axi_awlen        ,
		output wire [2 : 0]                        m00_axi_awsize       ,
		output wire [1 : 0]                        m00_axi_awburst      ,
		output wire                                m00_axi_awlock       ,
		output wire [3 : 0]                        m00_axi_awcache      ,
		output wire [2 : 0]                        m00_axi_awprot       ,
		output wire [3 : 0]                        m00_axi_awqos        ,
		output wire [C_M00_AXI_AWUSER_WIDTH-1 : 0] m00_axi_awuser       ,
		output wire                                m00_axi_awvalid      ,
		input wire                                 m00_axi_awready      ,
		output wire [C_M00_AXI_DATA_WIDTH-1 : 0]   m00_axi_wdata        ,
		output wire [C_M00_AXI_DATA_WIDTH/8-1 : 0] m00_axi_wstrb        ,
		output wire                                m00_axi_wlast        ,
		output wire [C_M00_AXI_WUSER_WIDTH-1 : 0]  m00_axi_wuser        ,
		output wire                                m00_axi_wvalid       ,
		input wire                                 m00_axi_wready       ,
		input wire [C_M00_AXI_ID_WIDTH-1 : 0]      m00_axi_bid          ,
		input wire [1 : 0]                         m00_axi_bresp        ,
		input wire [C_M00_AXI_BUSER_WIDTH-1 : 0]   m00_axi_buser        ,
		input wire                                 m00_axi_bvalid       ,
		output wire                                m00_axi_bready       ,
		output wire [C_M00_AXI_ID_WIDTH-1 : 0]     m00_axi_arid         ,
		output wire [C_M00_AXI_ADDR_WIDTH-1 : 0]   m00_axi_araddr       ,
		output wire [7 : 0]                        m00_axi_arlen        ,
		output wire [2 : 0]                        m00_axi_arsize       ,
		output wire [1 : 0]                        m00_axi_arburst      ,
		output wire                                m00_axi_arlock       ,
		output wire [3 : 0]                        m00_axi_arcache      ,
		output wire [2 : 0]                        m00_axi_arprot       ,
		output wire [3 : 0]                        m00_axi_arqos        ,
		output wire [C_M00_AXI_ARUSER_WIDTH-1 : 0] m00_axi_aruser       ,
		output wire                                m00_axi_arvalid      ,
		input wire                                 m00_axi_arready      ,
		input wire [C_M00_AXI_ID_WIDTH-1 : 0]      m00_axi_rid          ,
		input wire [C_M00_AXI_DATA_WIDTH-1 : 0]    m00_axi_rdata        ,
		input wire [1 : 0]                         m00_axi_rresp        ,
		input wire                                 m00_axi_rlast        ,
		input wire [C_M00_AXI_RUSER_WIDTH-1 : 0]   m00_axi_ruser        ,
		input wire                                 m00_axi_rvalid       ,
		output wire                                m00_axi_rready
	);
SYSTOLIC_ARRAY_v1_0_M00_AXI #
	(
		// Users to add parameters here
	.SYSTOLIC_SIZE     ( SYSTOLIC_SIZE     ),
	.DATA_WIDTH        ( DATA_WIDTH        ),
	.INOUT_WIDTH       ( INOUT_WIDTH       ),
	.IFM_RAM_SIZE      ( IFM_RAM_SIZE      ),
	.WGT_RAM_SIZE      ( WGT_RAM_SIZE      ),
	.OFM_RAM_SIZE_1    ( OFM_RAM_SIZE_1    ),
  .OFM_RAM_SIZE_2    ( OFM_RAM_SIZE_2    ),
	.MAX_WGT_FIFO_SIZE ( MAX_WGT_FIFO_SIZE ),
	.RELU_PARAM        ( RELU_PARAM        ),
  .Q                 ( Q                 ),
  .NUM_LAYER         ( NUM_LAYER         ),
  .ID_WIDTH          ( ID_WIDTH          ),
  .ADDR_WIDTH        ( ADDR_WIDTH        ),
  .LEN_WIDTH         ( LEN_WIDTH         ),


		// User parameters ends
		// Base address of targeted slave
		.C_M_TARGET_SLAVE_BASE_ADDR (C_M_TARGET_SLAVE_BASE_ADDR )  ,
		.C_M_AXI_BURST_LEN          (C_M_AXI_BURST_LEN          )  ,
		.C_M_AXI_ID_WIDTH           (C_M_AXI_ID_WIDTH           )  ,
		.C_M_AXI_ADDR_WIDTH         (C_M_AXI_ADDR_WIDTH         )  ,
		.C_M_AXI_DATA_WIDTH         (C_M_AXI_DATA_WIDTH         )  ,
		.C_M_AXI_AWUSER_WIDTH       (C_M_AXI_AWUSER_WIDTH       )  ,
		.C_M_AXI_ARUSER_WIDTH       (C_M_AXI_ARUSER_WIDTH       )  ,
		.C_M_AXI_WUSER_WIDTH        (C_M_AXI_WUSER_WIDTH        )  ,
		.C_M_AXI_RUSER_WIDTH        (C_M_AXI_RUSER_WIDTH        )  ,
		.C_M_AXI_BUSER_WIDTH        (C_M_AXI_BUSER_WIDTH        ) 
	) top_systolic
	(
//		input wire  INIT_AXI_TXN, // start transacsison
    .TXN_DONE      ( m00_axi_txn_done ) ,
    .ERROR         ( m00_axi_error    ) ,
    .M_AXI_ACLK    ( m00_axi_aclk     ) ,
    .M_AXI_ARESETN ( m00_axi_aresetn  ) ,
    .M_AXI_AWID    ( m00_axi_awid     ) ,
    .M_AXI_AWADDR  ( m00_axi_awaddr   ) ,
    .M_AXI_AWLEN   ( m00_axi_awlen    ) ,
    .M_AXI_AWSIZE  ( m00_axi_awsize   ) ,
    .M_AXI_AWBURST ( m00_axi_awburst  ) ,
    .M_AXI_AWLOCK  ( m00_axi_awlock   ) ,
    .M_AXI_AWCACHE ( m00_axi_awcache  ) ,
    .M_AXI_AWPROT  ( m00_axi_awprot   ) ,
    .M_AXI_AWQOS   ( m00_axi_awqos    ) ,
    .M_AXI_AWUSER  ( m00_axi_awuser   ) ,
    .M_AXI_AWVALID ( m00_axi_awvalid  ) ,
    .M_AXI_AWREADY ( m00_axi_awready  ) ,
    .M_AXI_WDATA   ( m00_axi_wdata    ) ,
    .M_AXI_WSTRB   ( m00_axi_wstrb    ) ,
    .M_AXI_WLAST   ( m00_axi_wlast    ) ,
    .M_AXI_WUSER   ( m00_axi_wuser    ) ,
    .M_AXI_WVALID  ( m00_axi_wvalid   ) ,
    .M_AXI_WREADY  ( m00_axi_wready   ) ,
    .M_AXI_BID     ( m00_axi_bid      ) ,
    .M_AXI_BRESP   ( m00_axi_bresp    ) ,
    .M_AXI_BUSER   ( m00_axi_buser    ) ,
    .M_AXI_BVALID  ( m00_axi_bvalid   ) ,
    .M_AXI_BREADY  ( m00_axi_bready   ) ,
    .M_AXI_ARID    ( m00_axi_arid     ) ,
    .M_AXI_ARADDR  ( m00_axi_araddr   ) ,
    .M_AXI_ARLEN   ( m00_axi_arlen    ) ,
    .M_AXI_ARSIZE  ( m00_axi_arsize   ) ,
    .M_AXI_ARBURST ( m00_axi_arburst  ) ,
    .M_AXI_ARLOCK  ( m00_axi_arlock   ) ,
    .M_AXI_ARCACHE ( m00_axi_arcache  ) ,
    .M_AXI_ARPROT  ( m00_axi_arprot   ) ,
    .M_AXI_ARQOS   ( m00_axi_arqos    ) ,
    .M_AXI_ARUSER  ( m00_axi_aruser   ) ,
    .M_AXI_ARVALID ( m00_axi_arvalid  ) ,
    .M_AXI_ARREADY ( m00_axi_arready  ) ,
    .M_AXI_RID     ( m00_axi_rid      ) ,
    .M_AXI_RDATA   ( m00_axi_rdata    ) ,
    .M_AXI_RRESP   ( m00_axi_rresp    ) ,
    .M_AXI_RLAST   ( m00_axi_rlast    ) ,
    .M_AXI_RUSER   ( m00_axi_ruser    ) ,
    .M_AXI_RVALID  ( m00_axi_rvalid   ) ,
    .M_AXI_RREADY  ( m00_axi_rready   ) ,
    .start_read    ( start_read       ) ,
    .done          ( done             )
	);
