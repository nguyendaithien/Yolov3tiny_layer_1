// generated case lines: address -> 256'bdata
module LUT #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 16
)(
	  input clk,
    input  [ADDR_WIDTH-1:0] address,
    output reg [DATA_WIDTH-1:0] data_out
);

  always @(posedge clk) begin
    case(address)
    32'd0 :  data_out = 256'b0000000001001001111100100000011100000011110110101111101111001100000010101100010100001011011110101111001100111010111100100101011011111100100111100000111001110101001010101010011111110001110011110000000111001101000000001011010111110110011101000000001100001111;
    32'd16 : data_out = 256'b0000000110011001111011000001011000000110110110111111101101111100000000000000010000010010100101101111110001110010000000110000100111110110011111000001111000010011000001011100011111101001101110110000001000000001000000011001011111111011111001110000011010111010;
    32'd32 : data_out = 256'b0000000011001110111101011001100100000100110010111111101011010100111101001011100000001011000101010000110001010110000101000011001100000010110000110000010000110111111001101100111111110010000100101111111111010100000000000101011000010001000101110000001110100010;
    32'd48 : data_out = 256'b1111110111110111000000110000100011111001100110111111101001000011000100100100000011111110111110101110110110011000111100111011110011111100101001111111111000001000000111100001000100000100011101100000010110000010000000011000010100000100010111010000100000001110;
    32'd64 : data_out = 256'b1111110101011111111111111010101111101011010000011111100001011101111110110011101000000000000011101111111100011101111001100000100111110001010110010000100001111000111110001111011011111111111011100000011001011011000000011100101000000001101101111111110001011001;
    32'd80 : data_out = 256'b0000000000111010111111111000000111101101000110111111101000110011111100000100111111111111110100000001001101011001001000000110000111111110000101011111001010010110111000100001100000000001011001000000001101010011000000001011101011111000011111101111100010011100;
    32'd96 : data_out = 256'b1111111110110100000011000100111000000010101000101111110111100111000011001000111111110101001100001111001011010001000001110000100000000001100011101111010000000001000011100011000000001101100101100000001101111000000000001000001100000110001011011111111111000010;
    32'd112 : data_out = 256'b1111110011011010000100111011000000001010010110111111100010101010111111110011011011101111111010010000010101010010111001011011010000000010000000111111001000001101111110011111010000010010001101010000010001011101000000010000101100000111111000011111001010000000;
    32'd128 : data_out = 256'b1111111001110000000010100101110100010001101000111111111000001101111101111000100111110011010111010000110010011000000011110011101011111111011001001110111111001101110111001100111100001010111100100000001011000000000000000001110111110111111001011111111000001101;
    32'd144 : data_out = 256'b1111110110011110111101010010010000000101001101010000001101100101000010111100101100001001101001001111010100001111111111011000001100000010110000000000100000111100111010101110000111110000100001001111111001100001000000001000000000000011000011010000001100001111;
    32'd160 : data_out = 256'b1111110100111110111011011100100100001010001010100000001111100011000000001000100100010010000101011111110111010111111111011000000111110111111111100001101010011011111110100011011011101001111101011111111001110111000000100010100011110011010001110000010100010011;
    32'd176 : data_out = 256'b1111101100100001111101110110100000000111101000010000000001111111111100111101100100001000010110010000101001011010000010110100000000000010101000000000000110100100000011000100110111110100101110100000000000110101000000010111111000010001000001100000000000000100;
    32'd192 : data_out = 256'b1111110001010110000001001001001011111001100111010000001001110101000100101100011011111110010101101110111010110100000001001110100011111111101100011111111001110111111110101000010000000010000011011111101101110101000000001111000111101110000110010000010001111100;
    32'd208 : data_out = 256'b1111101111001101000000000111010011101010010010110000000101111101111110111001010000000000001110101111111101001010111000010001111011110011111111010000110000011100111111111001000000000101010100101111101011111100000000011010010100001010001010011111101001000101;
    32'd224 : data_out = 256'b1111111001001011000000000100110011101010111010100000000101001111111011110100011000000000001110100001000101111011000100011100100111111111100110001111010000101111000100011101001000000001011110101111110110001100000000010100111111111010000011111111011100110000;
    32'd240 : data_out = 256'b1111110110110011000010000100101000000001011100010000001001000100000010011011111011110110100110011111010011110100000101110101010111111110001010111111010110100011111111111011010000001011010001111111110010101001000000001100010100010001011111000000000011011001;
    32'd256:  data_out = 256'b1111101110100001000100001111011000001001001011001111111101110001000000000000000011110000110100000000010101011001111010110000111000000010000000111111010100101111000000111101011100010011101110011111101111111000000000010101101111111110010001111111011010100010;
    32'd272:  data_out = 256'b1111110111111111000001101101000000001111110101000000000111101000111110000110000111110101101000110000100000110100111111111000111011111101100011001111000001001011000010101011011000001000101001101111110110100001000000001000010100000101110010110000000001011010;
    32'd288:  data_out = 256'b0000001110100111111101111100111100000100110111110000001010000111000001110010011000000101110100101111100101010110000001000000101100000001101011100000010101111010111001010100011011110111101011001111111111110100111111100100101000010001010011111111101101001001;
    32'd304:  data_out = 256'b0000010000101110111100110001100100000111001100000000010001100000000000100000100000001010100111010000000001100100111111110000001111111101010000100000110011100000111111000101011111101111111010011111111110100111111111101010010000001001001001011111111111111110;
    32'd320:  data_out = 256'b0000000000101000111110010011100000000101110010000000000111111100111101110110001100000100000101100000010111011000111111000101100100000011011010110000010011001111000010101011011011111001010000110000000000000110111111110100101111100110111100111111110111111000;
    32'd336:  data_out = 256'b0000010001010010000001000100011011111100110111010000001001001011000011001011100011111111100001001111010010010001000010101001001011111110101000011111110011001010111001001101001100000011011100001111111011111011111111000111010100000100011101110000000000000000;
    32'd352:  data_out = 256'b0000011000010111000000010001000111110010011001010000001010110100111111101000100000000001011101010000000100110010111100100111010011110101100101010000010000100111000000110111111000000011010100001111111010001010111110111000001000010011101101101111111111111100;
    32'd368:  data_out = 256'b0000010011101000000000000011011011110001110101100000010000000010111100110110110100000001001111110000101000011100111111010100011000000000011000101111110000001001000101011100011100000001011111001111111101000000111111001000001000001000010010111111111001001010;
    32'd384:  data_out = 256'b0000001100000100000001011110001000000000000000010000001001000101000001111100000011111001100000111111011011101111000100111001000011111111001100111111100111101000111100110100011100000110010011111111111110010110111111101111110111110101101010101111111110100101;
    32'd400:  data_out = 256'b0000010001111101000010111110100000000011010010010000000111011111000000010101111011110101110100000000010101110001111110111111010000000010101000101111100010000111000001111111011000001010111101001111111100111001111111101001111111110010000111011111110011011101;
    32'd416:  data_out = 256'b0000010000001001000001001101101100001001101001010000010000111011111110000000111011111001011100010000010011011100111101100011111011111100001000101111100111001011000110010111110100000110001110001111111101110111111111100000000100000100111000000000000100001110;
    32'd432 : data_out = 256'b1111111110100010000000000101101111111111111110000000000000000010111111111110101111111111111011111111111111101011000000000100110100000000000000000000000000000111000000000001001000000000001111010000000000110011111111111011000100000000000001000000000000000111;
   default: data_out = 256'd0;
endcase
end
endmodule
